package test_pkg;
 
 import uvm_pkg::*;

`include "uvm_macros.svh"

`include "trans.sv"
`include "seqs.sv"
`include "mon.sv"
`include "drv.sv"
`include "seqr.sv"


`include "agt.sv"
`include "scoreboard.sv"
`include "env.sv"

`include "base_test.sv"

endpackage