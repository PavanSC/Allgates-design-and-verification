interface intf(input bit clk);

  logic a;
  logic b;

  logic and_g;
  logic or_g;
  logic not_g;
  logic nor_g;
  logic nand_g;
  logic xor_g;
  logic xnor_g;


endinterface